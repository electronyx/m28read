`timescale 1ns / 1ps

//by M.Kachel
//
//BASED ON: https://github.com/sergachev/spi_mem_programmer
//The MIT License (MIT)
//
//Copyright (c) 2016 Ilia Sergachev

//Permission is hereby granted, free of charge, to any person obtaining a copy of this software and associated documentation files (the "Software"), to deal in the Software without restriction, including without limitation the rights to use, copy, modify, merge, publish, distribute, sublicense, and/or sell copies of the Software, and to permit persons to whom the Software is furnished to do so, subject to the following conditions:
//
//The above copyright notice and this permission notice shall be included in all copies or substantial portions of the Software.
//
//////////////////////////////////////////////////////////////////////////////////



//module spi_cmd(reset,SCLK,CS, SI_IO0,SO_IO1,WP_IO2,HOLD_IO3, 
//               busy,trigger, data_in_count,data_out_count,data_in,data_out,quad);
module spi_cmd(CLK,mem_clk,RST,CS, SI_IO0,SO_IO1,WP_IO2,HOLD_IO3, 
               busy,trigger, data_in_count,data_out_count,data_in,data_out,quad);
//
  input CLK;
  output  mem_clk;//serial clock
  input RST;
  //input SCLK; //serial clock - generated by PLL and also given to the output
  //input reset; //might be omitted  - same as power on
  output reg CS;
  inout SI_IO0; //serial input
  inout SO_IO1; //serial output
  inout WP_IO2; //write protect not used
  inout HOLD_IO3; //hold not used
  //all four IO0-3 are used for quad transfer
  
  output busy;
  
  input trigger;
  input [8:0] data_in_count; //into the memory - sending from FPGA
  input [3:0] data_out_count; //out of the memory  - received by FPGA
  input [79:0] data_in;
  output reg [47:0] data_out;
  input quad;
 
  wire [79:0]data_in_w;  
  assign   data_in_w=data_in;
  wire [3:0] DQ;

  reg [11:0] send_bit_cntr;
  reg [11:0] read_bit_cntr;
  
  wire [11:0] next_send_bit_cntr;
  assign next_send_bit_cntr=send_bit_cntr-1'b1;
  wire [11:0] next_read_bit_cntr;
  assign next_read_bit_cntr=read_bit_cntr-1'b1;
  
  
  //assign SI_IO0   = 
  reg OE; //output enable : 1-output, 0-input
  assign SI_IO0   =       OE?DQ[0]:1'bZ;
  assign SO_IO1   =       OE?DQ[1]:1'bZ;
  assign WP_IO2   =       OE?DQ[2]:1'bZ;
  assign HOLD_IO3 = quad?(OE?DQ[3]:1'bZ):1'b1; // has to be held 1 as 'hold' in non-quad mode
  
  
  wire [2:0] width = quad?3'b100:3'b001;
  //wire [2:0] width_1 = width -1'b1;


  parameter IDLE=4'b0000, SEND=4'b0001, READ=4'b0010, LAST_READ=4'b0011, WAIT_ONE_BEFORE_READ=4'b0100;
  reg [3:0] MEM_SPI_state;
  reg [3:0] next_MEM_SPI_state;
 
  reg [4:0] mem_clk_reg;
  
  assign mem_clk=mem_clk_reg[3];
  
  /*always@(posedge CLK) begin
     if(RST) mem_clk_reg<=4'b0011;
     else mem_clk_reg<={mem_clk_reg[2:0],mem_clk_reg[3]};
  end
*/

always@(posedge CLK) begin
   if(RST) begin
	   //mem_clk<=1'b0;
		CS<=1'b1;
		OE <= 1'b1;
		MEM_SPI_state<=IDLE;
	end
	else if(MEM_SPI_state==IDLE) begin
	  
		if(trigger && !busy ) begin
		   MEM_SPI_state<=SEND;
		   send_bit_cntr<=(data_in_count<<3)-1'b1;//load counter = bytes to bits
		   read_bit_cntr<=(data_out_count<<3)-1'b1;
			CS<=1'b0;
		end
      else begin
		  // mem_clk<=1'b0;
		   mem_clk_reg<=4'b0011;
		   CS<=1'b1;	
		   OE <= 1'b1;
		end
	end
	else if(MEM_SPI_state==SEND  ) begin
	   CS<=1'b0;
           if(mem_clk_reg==4'b0011) mem_clk_reg<=4'b0110;
		else if(mem_clk_reg==4'b0110) mem_clk_reg<=4'b1100;
		else if(mem_clk_reg==4'b1100) mem_clk_reg<=4'b1001;
		else if(mem_clk_reg==4'b1001) begin
		   mem_clk_reg<=4'b0011;
		   if(send_bit_cntr>width-1'b1) send_bit_cntr<=next_send_bit_cntr;
			else if(send_bit_cntr==12'h000 && data_out_count!=4'b0000) begin
			   MEM_SPI_state<=READ;
				OE<=1'b0;
			end
			else if(send_bit_cntr==12'h000 && data_out_count==4'b0000) MEM_SPI_state<=IDLE;
		end
		
   end
	else if(MEM_SPI_state==READ ) begin
	   CS<=1'b0;
		OE<=1'b0;
		
		     if(mem_clk_reg==4'b0011) mem_clk_reg<=4'b0110;
		else if(mem_clk_reg==4'b0110) mem_clk_reg<=4'b1100;
		else if(mem_clk_reg==4'b1100)  mem_clk_reg<=4'b1001;
		else if(mem_clk_reg==4'b1001) begin		
		   mem_clk_reg<=4'b0011;
	      if((read_bit_cntr>width-1'b1)) read_bit_cntr<=next_read_bit_cntr;
			else if(read_bit_cntr==(width-1'b1)) MEM_SPI_state<=IDLE;
			
			if(quad) data_out <= {data_out[43:0], SI_IO0, SO_IO1, WP_IO2, HOLD_IO3};
			else	   data_out <= {data_out[46:0], SO_IO1};
		   //mem_clk<=1'b1;
		end

	end


end

/*
//---------------------- CS handling
always@(posedge CLK) begin
   if(RST) CS=1'b1;
	else if(MEM_SPI_state==SEND || MEM_SPI_state==READ ||MEM_SPI_state==LAST_READ|| MEM_SPI_state==WAIT_ONE_BEFORE_READ ) CS=1'b0;
	else CS=1'b1;
end

//---------------------- send bit counter handling
always@(posedge CLK) begin
   if(RST) send_bit_cntr<=12'h000;
	else if(MEM_SPI_state == IDLE && trigger && !busy) send_bit_cntr<=(data_in_count<<3);//load counter = bytes to bits
   else if(SCK_fallingedge && MEM_SPI_state == SEND && (send_bit_cntr>width-1'b1) ) send_bit_cntr<=next_send_bit_cntr;
	
	

end
//---------------------- read bit counter handling
always@(posedge CLK) begin
   if(RST) read_bit_cntr<=12'h000;
	else if(MEM_SPI_state == IDLE && trigger && !busy) read_bit_cntr<=(data_out_count<<3);//load counter = bytes to bits
   else if(SCK_risingedge && MEM_SPI_state == READ && (read_bit_cntr>width-1'b1)) read_bit_cntr<=next_read_bit_cntr; //count 
end
*/
//---------------------- OE handling
//always@(posedge CLK) begin
//   if(RST) OE = 1'b1;
//	else if(MEM_SPI_state == READ ||MEM_SPI_state==LAST_READ ||MEM_SPI_state == WAIT_ONE_BEFORE_READ) OE = 1'b0;//??
//   else OE = 1'b1;
//end

assign busy = RST?1'b0:(MEM_SPI_state==SEND || MEM_SPI_state==READ ||MEM_SPI_state==LAST_READ|| MEM_SPI_state==WAIT_ONE_BEFORE_READ)?1'b1:1'b0;
////---------------------- busy handling
//always@(posedge CLK) begin
//   if(RST) busy=1'b0;
//	else if(MEM_SPI_state==SEND || MEM_SPI_state==READ ||MEM_SPI_state==LAST_READ|| MEM_SPI_state==WAIT_ONE_BEFORE_READ ) busy=1'b1;
//	else busy=1'b0;
//end



//----------------------SENDING DATA

wire [11:0] bitcntr3;
assign bitcntr3=send_bit_cntr-2'b11;
wire [11:0] bitcntr2;
assign bitcntr2=send_bit_cntr-2'b10;
wire [11:0] bitcntr1;
assign bitcntr1=send_bit_cntr-2'b01;


assign DQ[0] = quad?data_in_w[bitcntr3]: data_in_w[send_bit_cntr];
assign DQ[1] = quad?data_in_w[bitcntr2]: 1'bZ;
assign DQ[2] = quad?data_in_w[bitcntr1]: 1'bZ;
assign DQ[3] = quad?data_in_w[send_bit_cntr]:1'bZ;


//----------------------READING DATA
// always @(posedge CLK) begin
//	  if(RST)
//			data_out<=48'h000000000000;
//	  if(MEM_SPI_state==IDLE && trigger && !busy && SCK_fallingedge) data_out<=48'h000000000000;
//	  else if(SCK_fallingedge)
//         if(MEM_SPI_state==READ||MEM_SPI_state==LAST_READ) begin
//			  if(quad)
//				   data_out <= {data_out[43:0], SI_IO0, SO_IO1, WP_IO2, HOLD_IO3};
//				else
//				   data_out <= {data_out[46:0], SO_IO1};
//			end
// end


	 


endmodule
