`timescale 1ns / 1ps

//by M.Kachel
//
//BASED ON: https://github.com/sergachev/spi_mem_programmer
//The MIT License (MIT)
//
//Copyright (c) 2016 Ilia Sergachev

//Permission is hereby granted, free of charge, to any person obtaining a copy of this software and associated documentation files (the "Software"), to deal in the Software without restriction, including without limitation the rights to use, copy, modify, merge, publish, distribute, sublicense, and/or sell copies of the Software, and to permit persons to whom the Software is furnished to do so, subject to the following conditions:
//
//The above copyright notice and this permission notice shall be included in all copies or substantial portions of the Software.
//
//////////////////////////////////////////////////////////////////////////////////



//module spi_cmd(reset,SCLK,CS, SI_IO0,SO_IO1,WP_IO2,HOLD_IO3, 
//               busy,trigger, data_in_count,data_out_count,data_in,data_out,quad);
module spi_cmd(CLK,reset,SCLK,CS, SI_IO0,SO_IO1,WP_IO2,HOLD_IO3, 
               busy,trigger, data_in_count,data_out_count,data_in,data_out,quad);
//
  input CLK;
  input reset;
  input SCLK; //serial clock - generated by PLL and also given to the output
  //input reset; //might be omitted  - same as power on
  output reg CS;
  inout SI_IO0; //serial input
  inout SO_IO1; //serial output
  inout WP_IO2; //write protect not used
  inout HOLD_IO3; //hold not used
  //all four IO0-3 are used for quad transfer
  
  output reg busy;
  
  input trigger;
  input [8:0] data_in_count;
  input [3:0] data_out_count;
  input [260*8-1:0] data_in;
  output reg [47:0] data_out;
  input quad;
 
      
  reg [3:0] DQ = 4'b1111;

  reg [11:0] bit_cntr;
  reg [11:0] new_bit_cntr;
  wire [11:0] init_bit_cntr;
  assign init_bit_cntr=(data_in_count<<3)-1'b1;
  //assign SI_IO0   = 
  reg OE; //output enable : 1-output, 0-input
  assign SI_IO0   =       OE?DQ[0]:1'bZ;
  assign SO_IO1   =       OE?DQ[1]:1'bZ;
  assign WP_IO2   =       OE?DQ[2]:1'bZ;
  assign HOLD_IO3 = quad?(OE?DQ[3]:1'bZ):1'b1; // has to be held 1 as 'hold' in non-quad mode
  
 
  

  wire [2:0] width = 3'b001;//quad?4:1;



  parameter STATE_IDLE=4'b0000, STATE_SEND=4'b0001, STATE_READ=4'b0010,LAST_READ=4'b0011, STATE_WAIT_ONE_BEFORE_READ=4'b0100;
  reg [3:0] MEM_SPI_state;
  
  
  
  //reg [3:0] MEM_SPI_nextstate;
  //wire [11:0] init_bitcounter;
  //assign init_bitcounter=(data_in_count<<3)-1'b1;
  //init_bitcounter=data_in_count*8-1'b1;
  
  //start message
reg [2:0] SSELr; 
wire CSEL_FallingEdge = (SSELr[2:1]==2'b10); //message starts

//bit sampling on SCK falling edge
reg [2:0] SCKr;  
always @(posedge CLK) begin
   if(reset)begin
	   SCKr <= 3'b000;
      SSELr<= 3'b000;
	end
	else begin
	   SCKr <= {SCKr[1:0], SCLK};
      SSELr <= {SSELr[1:0], CS};
	end
end
wire SCK_risingedge =  (SCKr[2:1]==2'b01)?1:0;  // now we can detect SCK rising edges
wire SCK_fallingedge = (SCKr[2:1]==2'b10)?1:0;  // and falling edges
  
  //always @(posedge SCLK) begin
  always @(posedge CLK) begin
	  if(reset) begin
			MEM_SPI_state <= STATE_IDLE;
         OE   <= 1'b1;//lines as outputs
			busy <= 1'b1; //?
			CS   <=1'b1;
         bit_cntr <=12'h000;
	  end 
	  else begin
	     case(MEM_SPI_state)
				STATE_IDLE: begin
				OE <= 1'b1;
				   //trigger came but the controller is not yet busy -> go to send state
					if(trigger && !busy) begin
	
  //added if(SCK_fallingedge) - getting data out too soon?
                	if(SCK_fallingedge) begin 
						   MEM_SPI_state<=STATE_SEND; //you need to always send data first before reading
						   busy <= 1'b1;
						   bit_cntr <= init_bit_cntr;//(data_in_count<<3)-1'b1;
						end
						else begin
						   MEM_SPI_state<=MEM_SPI_state; //you need to always send data first before reading
						   busy <= busy;
						   bit_cntr <= bit_cntr;
						end
						
					end 
					else if(trigger && busy) //trigger came but controller busy
					begin
					   MEM_SPI_state<=STATE_IDLE;
						bit_cntr <= bit_cntr;
					end
					else if((!trigger&& busy) || (!trigger&& !busy)) //no trigger and controler busy - data transfer just finished			
					begin                                           //no trigger and controller not busy
						MEM_SPI_state<=STATE_IDLE;
						busy <= 1'b0;
						CS<=1'b1;
						bit_cntr <= bit_cntr;
					end	 
				end

				STATE_SEND: begin
				   CS<=1'b0;
					OE <= 1'b1;//OUTPUTS
					
					
					if(SCK_fallingedge) begin //if on the rising edge => timing problems come and sometimes data is 1bit delayed
					//if(SCK_risingedge) begin // rising edge SCK here is a falling edge of SCK in the MEMORY
					                         // so we prepare data here to be ready when the MEMORY will strobe
					
						/*if(quad) begin
							DQ[0] <= data_in[bit_cntr-2'b11];
							DQ[1] <= data_in[bit_cntr-2'b10];
							DQ[2] <= data_in[bit_cntr-2'b01];
							DQ[3] <= data_in[bit_cntr];
						end 
						else
							DQ[0] <= data_in[bit_cntr]; // 
					  */
					   //handle the bit counter
						if(bit_cntr>(width-1'b1)) begin // if the bitcounter is positive, send more data
							bit_cntr <= bit_cntr - width;
							MEM_SPI_state <= STATE_SEND;
						end				
						else if(bit_cntr==12'h000 && data_out_count!=4'b0000) begin //if bit counter became 0 and there is data to read
								 MEM_SPI_state <= STATE_WAIT_ONE_BEFORE_READ;                        //go to READ state
								 //MEM_SPI_state <= STATE_WAIT_ONE_BEFORE_READ;   
								 //OE <= 1'b0; //set to input -- NOT YET HERE, it will cause the last bit of SI to be 'Z'
				             //MEM_SPI_state <= STATE_READ;
								 bit_cntr <= (data_out_count<<3)-1'b1; 
								 //bit_cntr <= (data_out_count*8)-1'b1; 
						end
						else begin
								 MEM_SPI_state <= STATE_IDLE;
								 CS<=1'b1;
								 bit_cntr <= bit_cntr;
						end 
						
					end
					else begin
					   bit_cntr <= bit_cntr;
						MEM_SPI_state <= STATE_SEND;
				   end
				end
            STATE_WAIT_ONE_BEFORE_READ:begin
				   OE <= 1'b0; //set to input
					CS<=1'b0;
					bit_cntr <= bit_cntr;
					if(SCK_risingedge) MEM_SPI_state <= STATE_READ;
					else MEM_SPI_state <=STATE_WAIT_ONE_BEFORE_READ;
					
				
				end
				STATE_READ: begin
					OE <= 1'b0; //set to input
					CS<=1'b0;
					//if(SCK_fallingedge) begin
					if(SCK_risingedge) begin
					//
						if(bit_cntr>width-1'b1) begin
						   //CS<=1'b0;
							bit_cntr <= bit_cntr - width;
							MEM_SPI_state <= STATE_READ;
						end else begin
						   bit_cntr <= bit_cntr;
							MEM_SPI_state <= LAST_READ; //we still need to read on the next falling edge..
							//CS<=1'b0;//
						end
					end
					else begin
					   bit_cntr <= bit_cntr;
					   MEM_SPI_state <= STATE_READ;
					end
				end
            LAST_READ:
				begin
				   OE <= 1'b0; //set to input
				   CS<=1'b1;
					MEM_SPI_state <= STATE_IDLE;
					bit_cntr <= bit_cntr;
					if(SCK_risingedge) MEM_SPI_state <= STATE_IDLE;
					else  MEM_SPI_state <=LAST_READ;
				end
				default: begin
				   bit_cntr <= bit_cntr;
				   MEM_SPI_state <= STATE_IDLE;
               OE   <= 1'b1;//lines as outputs
			      CS   <=1'b1;
				end
			endcase
	  end
 end 
 
 wire [11:0] bitcntr3;
 assign bitcntr3=bit_cntr-2'b11;
 wire [11:0] bitcntr2;
 assign bitcntr2=bit_cntr-2'b10;
 wire [11:0] bitcntr1;
 assign bitcntr1=bit_cntr-2'b01;

 
 always@(posedge SCLK) begin
	 if(MEM_SPI_state==STATE_SEND)
	 begin 
		if(quad) begin
			DQ[0] <= data_in[bitcntr3];
			DQ[1] <= data_in[bitcntr2];
			DQ[2] <= data_in[bitcntr1];
			DQ[3] <= data_in[bit_cntr];
		end 
		else
			DQ[0] <= data_in[bit_cntr]; // 
	 end
 end

 always @(negedge SCLK or posedge reset) begin
	  if(reset)
			data_out<=48'h000000000000;
	  else
			//if(MEM_SPI_state==STATE_READ|| MEM_SPI_state==LAST_READ ) begin
         if(MEM_SPI_state==STATE_READ || MEM_SPI_state==LAST_READ ) begin
			  			  
			  if(quad)
				   data_out <= {data_out[43:0], SI_IO0, SO_IO1, WP_IO2, HOLD_IO3};
				else
				   data_out <= {data_out[46:0], SO_IO1};
			end
			//else if(MEM_SPI_state==STATE_WAIT_ONE_BEFORE_READ) data_out<=48'h000000000000;
 end

	 


endmodule
